BAT_MaxDisChgCurr , Bat.BusCurr, float
DC_FailSt_Inverted , Bat.BusVolt, float
