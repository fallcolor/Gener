TM_InvTemp, TM.InvTemp, int16_T
BAT_Volt, Bat.BusVolt, float
TM_EnergyActl, TM.EneAct
VCU_SpdSet, Set.vehSpd, float
TM_Volt_C, TM.VoltC, float
TM_Efficency, TM.Eff, float
TM_CtrlMode, TM.CM, avd